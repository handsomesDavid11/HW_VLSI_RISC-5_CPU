module ALU_ctrl(
     




);



endmodule